library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity template is
	port(
		Buttons : in std_logic_vector(3 downto 0);  -- Button 3 to Button 0
	Switches : in std_logic_vector(7 downto 0); -- Switch 7 to switch 0
		Clock50, Clock14 : in std_logic;  -- both clocks
		LED_A : out std_logic_vector(7 downto 0);  -- From LED 7 to LED 0
		LED_B : out std_logic_vector(7 downto 0);  -- From LED 7 to LED 0
		Segment1, Segment2, Segment3, Segment4 : out	std_logic_vector(7 downto 0)  -- From DP (7) to A (0) as defined in the docs 
		-- The pinheader needs to be defined by the user
	);
end entity;

architecture arch of template is

begin
	-- Place your architecture code here ...
end architecture;
